interface intf(input logic clk,rst);
logic mod;
logic clk;
logic rst;
logic[2:0] count;
endinterface

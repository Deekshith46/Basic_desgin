interface intf();
bit clk,rst;
logic mod;
logic[2:0] count;
endinterface

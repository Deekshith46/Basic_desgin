module test;
reg   [31:0]   instruction; // 32-bit instruction [1:0]
wire [1:0] bc_o; // bit class
wire        ct_o; //class type
wire [4:0]   opcode_o; //opcod
wire [4:0]   rd_addr;
wire [4:0]   rs1_addr;
wire [4:0]   rs2_addr;
wire [13:0]  immediate;
wire [18:0]  jump_imm;
wire [23:0]  system_op;


decoder dut(.instruction(instruction),
            .bc_o(bc_o),
            .ct_o(ct_o),
            .opcode_o(opcode_o),
            .rs1_addr(rs1_addr),
            .rs2_addr(rs2_addr),
            .rd_addr(rd_addr),
            .immediate(immediate),
            .jump_imm(jump_imm),
            .system_op(system_op));

        initial begin
            $shm_open("decoder.shm");
            $shm_probe("ACTMF");
        end

        initial begin
            instruction = 32'b00_0_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b00_0_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b00_0_00010_00011_00001_00010_0000_00000;//SUB
              #10
               instruction = 32'b00_0_00011_11010_00001_00010_0000_00000;//MUL
#10
                instruction = 32'b00_0_00100_11010_00001_00010_0000_00000;//SMUIL
#10
                 instruction = 32'b00_0_00101_00011_00001_00010_0000_00000;//DIV
#10
                  instruction = 32'b00_0_00110_00011_00001_00010_0000_00000;//IDIV
#10
                   instruction = 32'b00_0_00111_00011_00001_00010_0000_00000;//AND
#10
                    instruction = 32'b00_0_01000_00011_00001_00010_0000_00000;//OR

//////////////////////////////////I_TYPE//////////////////////////////////////////////////
            instruction = 32'b00_1_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b00_1_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b00_1_00010_00011_00001_00010_0000_00000;//SUB
              #10
               instruction = 32'b00_1_00011_11010_00001_00010_0000_00000;//MUL
#10
                instruction = 32'b00_1_00100_11010_00001_00010_0000_00000;//SMUIL
#10
                 instruction = 32'b00_1_00101_00011_00001_00010_0000_00000;//DIV
#10
                  instruction = 32'b00_1_00110_00011_00001_00010_0000_00000;//IDIV
#10
                   instruction = 32'b00_1_00111_00011_00001_00010_0000_00000;//AND
#10
                    instruction = 32'b00_1_01000_00011_00001_00010_0000_00000;//OR

///////////////////////////////////////////////LOAD_TYPE/////////////////////////////////////////
 instruction = 32'b01_0_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b01_0_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b01_0_00010_00011_00001_00010_0000_00000;//SUB
              #10
               instruction = 32'b01_0_00011_11010_00001_00010_0000_00000;//MUL
#1
                instruction = 32'b01_0_00100_11010_00001_00010_0000_00000;//SMUIL
#10
                 instruction = 32'b01_0_00101_00011_00001_00010_0000_00000;//DIV
#10
                  instruction = 32'b01_0_00110_00011_00001_00010_0000_00000;//IDIV
#10
                   instruction = 32'b01_0_00111_00011_00001_00010_0000_00000;//AND
#10
                    instruction = 32'b01_0_01000_00011_00001_00010_0000_00000;//OR
///////////////////////////////////////STORE_TYPE////////////////////////////////////////////////////////////////////////
instruction = 32'b01_1_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b01_1_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b01_1_00010_00011_00001_00010_0000_00000;//SUB
              #10
               instruction = 32'b01_1_00011_11010_00001_00010_0000_00000;//MUL
#1
                instruction = 32'b01_1_00100_11010_00001_00010_0000_00000;//SMUIL
#10
                 instruction = 32'b01_1_00101_00011_00001_00010_0000_00000;//DIV
#10
                  instruction = 32'b01_1_00110_00011_00001_00010_0000_00000;//IDIV
#10
                   instruction = 32'b01_1_00111_00011_00001_00010_0000_00000;//AND
#10
                    instruction = 32'b01_1_01000_00011_00001_00010_0000_00000;//OR
////////////////////////////////////////////BRANCH/////////////////////////////////////////////////////////////////
instruction = 32'b10_0_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b10_0_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b10_0_00010_00011_00001_00010_0000_00000;//SUB
              #10
               instruction = 32'b10_0_00011_11010_00001_00010_0000_00000;//MUL
#1
                instruction = 32'b10_0_00100_11010_00001_00010_0000_00000;//SMUIL
#10
                 instruction = 32'b10_0_00101_00011_00001_00010_0000_00000;//DIV
#10
                  instruction = 32'b10_0_00110_00011_00001_00010_0000_00000;//IDIV
#10
                   instruction = 32'b10_0_00111_00011_00001_00010_0000_00000;//AND
#10
                    instruction = 32'b10_0_01000_00011_00001_00010_0000_00000;//OR
///////////////////////////////////////////////JUMP////////////////////
instruction = 32'b10_1_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b10_1_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b10_1_00010_00011_00001_00010_0000_00000;//SUB
              #10

             instruction = 32'b10_1_00011_11010_00001_00010_0000_00000;//MUL
//////////////////////////////////SYSTEM_OPERATION/////////////////
instruction = 32'b11_0_00000_00011_00001_00010_0000_00000;//ADD
#10
             instruction = 32'b11_0_00001_00011_00001_00010_0000_00000;//ADDU
             #10

              instruction = 32'b11_0_00010_00011_00001_00010_0000_00000;//SUB
              #10
instruction = 32'b11_0_00011_11010_00001_00010_0000_00000;
#200
             $finish();
        end

endmodule   

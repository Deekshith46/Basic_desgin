interface intf(input logic clk,rst);
logic mod;
logic[2:0] count;
endinterface
